$display("Hello World");
$display("New");
$`timescale 1ps/1ps